module smart_traffic(
    input clk,
    input reset,
    input pedestrian,
    input ambulance,
    input [1:0] traffic_density,
    output reg red,
    output reg yellow,
    output reg green
);

reg [3:0] state;
reg [7:0] counter;

parameter RED=0, GREEN=1, YELLOW=2, PEDESTRIAN=3, AMBULANCE=4;

always @(posedge clk or posedge reset)
begin
    if(reset)
    begin
        state <= RED;
        counter <= 0;
    end
    else
    begin
        counter <= counter + 1;

        case(state)

        RED:
        begin
            if(ambulance) state <= AMBULANCE;
            else if(counter==5) begin state<=GREEN; counter<=0; end
        end

        GREEN:
        begin
            if(ambulance) state <= AMBULANCE;
            else if(pedestrian) state <= PEDESTRIAN;
            else if(counter == (traffic_density==2'b11 ? 15:8))
            begin
                state <= YELLOW;
                counter<=0;
            end
        end

        YELLOW:
        begin
            if(counter==3) begin state<=RED; counter<=0; end
        end

        PEDESTRIAN:
        begin
            if(counter==6) begin state<=RED; counter<=0; end
        end

        AMBULANCE:
        begin
            if(counter==10) begin state<=RED; counter<=0; end
        end

        endcase
    end
end

always @(*)
begin
    red=0; yellow=0; green=0;

    case(state)
    RED: red=1;
    GREEN: green=1;
    YELLOW: yellow=1;
    PEDESTRIAN: red=1;
    AMBULANCE: green=1;
    endcase
end

endmodule